module mux_2_to_1_v2 (
   input      a
  ,input      b
  ,input      sel
  ,output reg y
);

  always_comb
    if(sel)
      y = b;
    else
      y = a;
  
endmodule

// -------------------------------------------------------------------------- //
// Corresponding ciruit:
// -------------------- 
//  
//      |\
//  a --| \
//      |  |
//      |  |-- y
//      |  |
//  b --| /
//      |/
//
// -------------------------------------------------------------------------- //

