module mux_16_to_1 (
   input      [15:0] i
  ,input       [3:0] sel
  ,output reg        y
);

  always_comb
    case(sel)
      4'h0: y = i[ 0];
      4'h1: y = i[ 1];
      4'h2: y = i[ 2];
      4'h3: y = i[ 3];
      4'h4: y = i[ 4];
      4'h5: y = i[ 5];
      4'h6: y = i[ 6];
      4'h7: y = i[ 7];
      4'h8: y = i[ 8];
      4'h9: y = i[ 9];
      4'hA: y = i[10];
      4'hB: y = i[11];
      4'hC: y = i[12];
      4'hD: y = i[13];
      4'hE: y = i[14];
      4'hF: y = i[15];
    endcase
    
endmodule


// -------------------------------------------------------------------------- //
// Corresponding ciruit:
// -------------------- 
//  
//          |\
//  i[ 0] --| \
//          |  |
//  i[ 1] --|  |
//          |  |
//  i[ 2] --|  |
//          |  |
//  i[ 3] --|  |
//          |  |
//  i[ 4] --|  |
//          |  |
//  i[ 5] --|  |
//          |  |
//  i[ 6] --|  |
//          |  |
//  i[ 7] --|  |
//          |  |-- y
//  i[ 8] --|  |
//          |  |
//  i[ 9] --|  |
//          |  |
//  i[10] --|  |
//          |  |
//  i[11] --|  |
//          |  |
//  i[12] --|  |
//          |  |
//  i[13] --|  |
//          |  |
//  i[14] --|  |
//          |  |
//  i[15] --| /
//          |/
//
// -------------------------------------------------------------------------- //